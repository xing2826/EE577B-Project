// This is input channel for Clock Wise, which contains 2 virtual channel (input buffer)
`include "./ channelbuffer/ Input_ChannelBuffer.v"

module CW_Input_Channel (
    ports
);
    
endmodule