

module NIC (
    ports
);
    
endmodule