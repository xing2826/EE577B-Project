//the module shown in ''2022fall_cardinal_router.pdf' figure 3 
//containing 4 RTR and 2 PER modules.

module gold_router (
    input cwsi,
    input [63:0]cwdi,
    input ccwsi,
    input [63:0]ccwdi,
    input pesi,
    input pedi[63:0],
    input cwro,
    input ccwro,
    input pero,
    output cwri,
    output ccwri,
    output peri,
    output cwso,
    output [63:0]cwdo,
    output ccwso,
    output [63:0]ccwdo,
    output peso,
    output [63:0]pedo
);
    
endmodule