//the ring structual of the router, consisted by 4 gold_router modules. 
//the ring connnects to 4 processors so that they can communicate through the ring router.

module gold_ring (
    ports
);
    
endmodule