// The input and output PE channel use the same structual
//hence only one module designed below and instantiate 2 time in gold_router.v

module PER (
    ports
);
    
endmodule