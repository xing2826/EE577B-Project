// The CW and CCW in/out channel use the same structual
//hence only one module designed below and instantiate 4 time in gold_router.v

module RTR (
    ports
);
    
endmodule